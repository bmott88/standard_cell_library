** sch_path: /home/bmott/standard_cell_library/xsch/ip/inv/inv.sch
.subckt inv in out VDD VSS
*.ipin in
*.opin out
*.iopin VDD
*.iopin VSS
XMN out in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XMP out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
**.ends
.end
