** sch_path: /home/bmott/standard_cell_library/xsch/ip/tgate/tgate_6t.sch
**.subckt tgate_6t VDD VSS a b en
*.iopin a
*.iopin b
*.ipin en
*.iopin VDD
*.iopin VSS
x1 en selb VDD VSS inv
x2 selb sel VDD VSS inv
x3 a b sel selb VDD VSS tgate_2t
**.ends

* expanding   symbol:  ip/inv/inv.sym # of pins=4
** sym_path: /home/bmott/standard_cell_library/xsch/ip/inv/inv.sym
** sch_path: /home/bmott/standard_cell_library/xsch/ip/inv/inv.sch
.subckt inv in out VDD VSS
*.ipin in
*.opin out
*.iopin VDD
*.iopin VSS
XMN out in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XMP out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0
+ mult=1 m=1
.ends


* expanding   symbol:  ip/tgate/tgate_2t.sym # of pins=6
** sym_path: /home/bmott/standard_cell_library/xsch/ip/tgate/tgate_2t.sym
** sch_path: /home/bmott/standard_cell_library/xsch/ip/tgate/tgate_2t.sch
.subckt tgate_2t a b sel selb VDD VSS
*.iopin a
*.iopin b
*.iopin VDD
*.iopin VSS
*.ipin sel
*.ipin selb
XMP a selb b VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad=0.58 as=0.58 pd=4.58 ps=4.58 nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0 mult=1
+ m=1
XMN a sel b VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
.ends

.end
