* NGSPICE file created from tgate_2t.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_E5WSWT B D S G
X0 S G D B sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_EUN5X2 B D S G
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt tgate_2t a b sel selb VDD VSS
XXMN VSS a b sel sky130_fd_pr__nfet_01v8_E5WSWT
XXMP VDD a b selb sky130_fd_pr__pfet_01v8_EUN5X2
.ends

