magic
tech sky130A
magscale 1 2
timestamp 1766075075
<< viali >>
rect -290 1246 -8 1280
rect -290 -106 -8 -72
<< metal1 >>
rect -360 1280 62 1316
rect -360 1246 -290 1280
rect -8 1246 62 1280
rect -360 1216 62 1246
rect -290 1086 -244 1216
rect -192 1138 -106 1184
rect -290 1036 -176 1086
rect -210 708 -176 1036
rect -122 758 -88 1086
rect -122 708 -8 758
rect -182 306 -116 650
rect -54 256 -8 708
rect -210 130 -176 256
rect -290 80 -176 130
rect -122 206 -8 256
rect -122 80 -88 206
rect -290 -42 -244 80
rect -192 -10 -106 36
rect -360 -72 62 -42
rect -360 -106 -290 -72
rect -8 -106 62 -72
rect -360 -142 62 -106
use sky130_fd_pr__nfet_01v8_E5WSWT  XMN
timestamp 1766075075
transform 1 0 -149 0 1 168
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_ELW5X2  XMP
timestamp 1766074289
transform 1 0 -149 0 1 897
box -211 -419 211 419
<< labels >>
rlabel metal1 -182 306 -116 650 1 in
port 0 n
rlabel metal1 -54 206 -8 758 1 out
port 1 n
rlabel metal1 -360 1280 62 1316 1 VDD
port 2 n
rlabel metal1 -360 -142 62 -106 1 VSS
port 3 n
<< end >>
