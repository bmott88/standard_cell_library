magic
tech sky130A
timestamp 1766176949
<< metal1 >>
rect -1 679 632 729
rect -1 0 632 50
use inv  inv_0 ~/standard_cell_library/mag/inv
timestamp 1766075075
transform 1 0 179 0 1 71
box -180 -71 31 658
use inv  inv_1
timestamp 1766075075
transform 1 0 390 0 1 71
box -180 -71 31 658
use tgate_2t  tgate_2t_0 ~/standard_cell_library/mag/tgate_2t
timestamp 1766176949
transform 1 0 443 0 1 348
box -22 -348 189 381
<< end >>
