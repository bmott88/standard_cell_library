* NGSPICE file created from inv.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_E5WSWT B D S G
X0 S G D B sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_ELW5X2 B D S G
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt inv in out VDD VSS
XXMN VSS VSS out in sky130_fd_pr__nfet_01v8_E5WSWT
XXMP VDD VDD out in sky130_fd_pr__pfet_01v8_ELW5X2
.ends

