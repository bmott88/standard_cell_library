** sch_path: /home/bmott/tt_relative_path_test/xsch/tb/inv/inv_tb.sch
**.subckt inv_tb
x1 net1 in out GND inv
* noconn out
V1 in GND 1.8
V2 net1 GND 1.8
**** begin user architecture code
.lib /opt/pdk/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.control
set wr_singlescale
set wr_vecnames

dc V1 0 1.8 1m
wrdata OUTPUT.csv v(out)
quit
.endc


**** end user architecture code
**.ends

* expanding   symbol:  ip/inv/inv.sym # of pins=4
** sym_path: /home/bmott/tt_relative_path_test/xsch/ip/inv/inv.sym
** sch_path: /home/bmott/tt_relative_path_test/xsch/ip/inv/inv.sch
.subckt inv VDD in out VSS
*.ipin in
*.opin out
*.iopin VDD
*.iopin VSS
XM2 out in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM11 out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
.ends

.GLOBAL GND
.end
